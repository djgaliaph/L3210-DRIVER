��[ M a i n ]  
 C a p t i o n 	 = " I n s t a l l   N a v i   [ % P R O D U C T _ N A M E % ] "  
 B T N _ N e x t 	 = " N � s t a "  
  
 ; �% 
 B T N _ N e x t S t e p 	 	 = " N � s t a "  
 B T N _ S t a r t S e t t i n g 	 = " N � s t a "  
 B T N _ S t a r t 	 	 = " N � s t a "  
 B T N _ R e t r y   	 	 = " F � r s � k   i g e n "  
 B T N _ A b o r t 	 	 = " H o p p a   � v e r "  
 B T N _ R e c h e c k 	 	 = " B e k r � f t a   i g e n "  
 B T N _ A c c e p t 	 	 = " A c c e p t e r a "  
 B T N _ E x i t 	 	 = " A v s l u t a "  
 B T N _ A g r e e 	 	 = " G o d k � n n e r "  
  
 B T N _ B a c k 	 = " B a k � t "  
 B T N _ I n s t a l l 	 = " I n s t a l l e r a "  
 B T N _ C a n c e l 	 = " A v b r y t "  
 B T N _ F i n i s h 	 = " S l u t f � r "  
 B T N _ S k i p 	 = " H o p p a   � v e r "  
 B T N _ A p p l y 	 = " V e r k s t � l l "  
 B T N _ R e g i s t 	 = " R e g i s t r e r a "  
 B T N _ R e s t a r t 	 = " M o d e l l � t e r s t � l l n i n g "  
 B T N _ N W D i a g             = " D e t a l j e r "  
 B T N _ R e n e w a l   	 = " U p p d a t e r a "  
 B T N _ Y e s                   = " N � s t a "  
 B T N _ N o                     = " S t � n g "  
 P D M _ L a n g u a g e 	 = " S p r � k "  
 P D M _ S u p p o r t 	 = " S u p p o r t "  
 D L G _ C a n c e l 	 = " � r   d u   s � k e r   p �   a t t   d u   v i l l   a v b r y t a ? "  
 L B L _ W i f i 	 = " A n s l u t   v i a   t r � d l � s t   n � t v e r k   ( W i - F i ) "  
 L B L _ R e c o m m e n d e d 	 = " ( r e k o m m e n d e r a s ) "  
  
 L B L _ E n v C h e c k         = " K o n t r o l l e r a r   m i l j � n . . . "    
 L B L _ D e l D e v M e s s a g e     = " K o n t r o l l e r a r   m i l j � n . . . "    
 L B L _ D e l D e v C a u t i o n   =   " K o n t r o l l e n   k a n   t a   t i d .   R � r   i n t e   s k r i v a r e n   o c h   d a t o r n . "    
 L B L _ D e l D e v C a u t i o n   =   " "  
 L B L _ R e s t a r t 	 = " D u   m � s t e   s t a r t a   o m   d a t o r n   f � r   a t t   a n v � n d a   p r o g r a m m e t . "  
  
 [ F o r M a c ]  
 T I T L E 	 = " L � g g   t i l l   s k r i v a r e "  
 O p t i o n C b x 	 = " L a d d a   n e r   d e n   s e n a s t e   p r o g r a m v a r a n   f r � n   E p s o n "  
 ; O p t i o n C b x E x p 	 = " A k t i v e r a   i n s t a l l a t i o n   o c h   u p p d a t e r i n g   a v   p r o g r a m v a r a   s o m   d u   k a n   a n v � n d a . "  
 Q _ E x i s t M s g 	 = " F � r   n � r v a r a n d e   � r   A i r P r i n t - d r i v r u t i n e n   v a l d .   D u   k a n   a n v � n d a   v � r   p r o d u k t s   a l l a   f u n k t i o n e r   o m   d u   i   s t � l l e t   v � l j e r   E p s o n - d r i v r u t i n e n   g e n o m   a t t   k l i c k a   p �   k n a p p e n   h � r   n e d a n f � r . "  
 Q _ E x i s t A P B t n 	 = " A i r P r i n t "  
 Q _ E x i s t E P B t n 	 = " E p s o n "  
 Q _ N o E x i s t M s g 	 = " K l i c k a   p �   [ O K ]   f � r   a t t   l � g g a   t i l l   E p s o n   u t s k r i f t s k �   t i l l   u t s k r i f t s l i s t a n . "  
 Q _ N o E x i s t B t n 	 = " O K "  
 Q _ F a i l u r e M s g 	 = " R e g i s t r e r i n g   a v   s k r i v a r e   m i s s l y c k a d e s .   K l i c k a   p �   O K   o c h   r e g i s t r e r a   s e d a n   s k r i v a r e n   i g e n . "  
 Q _ F a i l u r e B t n 	 = " O K "  
 T e s t _ F a i l u r e M s g 	 = " T e s t u t s k r i f t   m i s s l y c k a d e s .   R e g i s t r e r a   s k r i v a r e n   i g e n . "  
 Q _ P r i n t e r N o t F o u n d   = " S k r i v a r e n   h i t t a d e s   i n t e . "  
  
 [ L e f t P r o g r e s s ]  
 S T R _ E u r a 	 = " L i c e n s a v t a l "  
 S T R _ S y s t e m C h e c k 	 = " V � l j   a l t e r n a t i v "  
 S T R _ I n s t a l l 	 = " I n s t a l l a t i o n "  
 S T R _ C o n n e c t i o n 	 = " I n s t a l l a t i o n "  
 S T R _ A d d I n s t a l l 	 = " K o m p l e t t e r a n d e   i n s t a l l a t i o n "    
 S T R _ F i n i s h 	 = " S l u t f � r "  
 ; �% 
 S T R _ O p e C h e c k 	 = " K o n t r o l l e r a   f u n k t i o n e r "  
  
 ; �% 
 [ e R e g _ A ]  
 P A T H E X E _ W 	 = " \ A p p s \ R e g i s t e r \ e R e g L a u n c h e r . e x e "  
 P A R A M _ W 	 	 = " / L a n g : U S "  
 P A T H E X E _ M 	 = " / A p p s / R e g i s t e r / E p s o n R e g R e d i r e c t . a p p "  
  
 [ S u p p o r t L i n k _ A ]  
 P A T H E X E _ M 	 = " / A p p s / S u p p o r t L i n k / U S / G u i d e . p k g "  
  
 [ S t a r t M e n u ]  
 T I T L E 	 = " I n s t a l l   N a v i "  
 L N K _ S t a r t 	 = " S t a r t   o c h   a n s l u t n i n g "  
 H L P _ S t a r t 	 = " K l i c k a   h � r   n � r   d u   v i l l   s t a r t a   i n s t a l l a t i o n s p r o c e s s e n ,   i n s t a l l e r a   p r o g r a m v a r a n   o c h   k o n f i g u r e r a   n � t v e r k s i n s t � l l n i n g a r . "  
 L N K _ G u i d e 	 = " E n d a s t   f � r   s y s t e m a d m i n i s t r a t � r e r "  
 H L P _ G u i d e 	 = " K l i c k a   h � r   o m   d u   v i l l   v i s a   s k r i v a r e n s   h a n d b o k   o m   m a s k i n v a r u i n s t a l l a t i o n   ( P D F )   o c h   a n d r a   a d m i n i s t r a t i v a   i n s t � l l n i n g a r . "  
 L N K _ M a n u a l 	 = " I n f o r m a t i o n   f � r   h a n d b � c k e r   o c h   p r o g r a m "  
 H L P _ M a n u a l 	 = " K l i c k a   h � r   f � r   a t t   f �   i n f o r m a t i o n   o m   h a n d b � c k e r ,   d e   v a n l i g a s t e   p r o g r a m m e n   s � s o m   s k r i v a r d r i v r u t i n e r   o c h   s � k v � g a r   t i l l   d e s s a   p r o g r a m   s o m   f i n n s   p �   p r o g r a m v a r a n s   c d - s k i v a   s �   a t t   d u   k a n   i n s t a l l e r a   d e m   m a n u e l l t . "  
  
 [ A s s i s t a n t ]  
 A S S _ N o C o n n e c t _ F u l l 	 = " < I n f o r m a t i o n > \ n D e t   f i n n s   U S B - k a b e l a n s l u t n i n g   f � r   a t t   a n s l u t a   p r o d u k t e n   o c h   d a t o r n . "  
 A S S _ N o N e t w o r k _ F u l l 	 = " < I n f o r m a t i o n > \ n D e t   f i n n s   t r � d l � s   L A N - a n s l u t n i n g   ( W i - F i )   f � r   a t t   a n s l u t a   p r o d u k t e n   o c h   d a t o r n . "  
 A S S _ N o W i F i _ F u l l 	 	 = " < I n f o r m a t i o n > \ n D u   k a n   a n s l u t a   p r o d u k t e n   o c h   d a t o r n   d i r e k t . "  
 A S S _ N o W A C _ F u l l 	 	 = " < I n f o r m a t i o n > \ n D u   k a n   a n s l u t a   p r o d u k t e n   o c h   d a t o r n   v i a   n � t v e r k . "  
 A S S _ O k W A C _ F u l l 	 	 = " < I n f o r m a t i o n > \ n D u   k a n   a n s l u t a   p r o d u k t e n   o c h   d a t o r n   v i a   t r � d l � s t   L A N   ( W i - F i ) . "  
  
 A S S _ N o C o n n e c t _ O n l y W i F i 	 = " < I n f o r m a t i o n > \ n D e t   f i n n s   U S B - k a b e l a n s l u t n i n g   f � r   a t t   a n s l u t a   p r o d u k t e n   o c h   d a t o r n . "  
 A S S _ N o N e t w o r k _ O n l y W i F i 	 = " < I n f o r m a t i o n > \ n D e t   f i n n s   t r � d l � s   L A N - a n s l u t n i n g   ( W i - F i )   f � r   a t t   a n s l u t a   p r o d u k t e n   o c h   d a t o r n . "  
 A S S _ N o W i F i _ O n l y W i F i 	 = " < I n f o r m a t i o n > \ n D u   k a n   a n s l u t a   p r o d u k t e n   o c h   d a t o r n   d i r e k t . "  
 A S S _ N o W A C _ O n l y W i F i 	 = " < I n f o r m a t i o n > \ n D u   k a n   a n s l u t a   p r o d u k t e n   o c h   d a t o r n   v i a   n � t v e r k . "  
 A S S _ O k W A C _ O n l y W i F i 	 = " < I n f o r m a t i o n > \ n D u   k a n   a n s l u t a   p r o d u k t e n   o c h   d a t o r n   v i a   t r � d l � s t   L A N   ( W i - F i ) . "  
 A S S _ N o W i F i _ A l e r t 	 = " D a t o r n   � r   i n t e   a n s l u t e n   t i l l   n � g o t   n � t v e r k .   A n s l u t   d a t o r n   t i l l   e t t   n � t v e r k   f � r   a t t   s k r i v a   u t   e l l e r   s k a n n a   ( i   f � r e k o m m a n d e   f a l l )   � v e r   n � t v e r k e t . "  
 A S S _ O n l y W i F i _ A l e r t 	 = " D a t o r n   � r   a n s l u t e n   t i l l   e t t   W i - F i   D i r e c t - n � t v e r k .   D u   k a n   a n v � n d a   e n   U S B -   e l l e r   W i - F i   D i r e c t - a n s l u t n i n g   f � r   a t t   s k r i v a   u t   e l l e r   s k a n n a   ( i   f � r e k o m m a n d e   f a l l ) . "  
  
 [ S e l e c t M o d e l ]  
 T I T L E = " V � l j   d i n   p r o d u k t "  
 T X T _ B o d y = " V � l j   d i n   p r o d u k t   f r � n   l i s t a n . "  
  
 [ F o r A d m i n ]  
 T I T L E 	 = " E n d a s t   f � r   s y s t e m a d m i n i s t r a t � r e r "  
 S U B _ T i t l e 	 = " "  
 B T N _ H S G 	 = " H a n d b o k   f � r   m a s k i n v a r u i n s t a l l a t i o n "  
  
 [ V i e w M a n u a l ]  
 T I T L E 	 = " I n f o r m a t i o n   f � r   h a n d b � c k e r   o c h   p r o g r a m "  
 S U B _ T i t l e 	 = " "  
 B T N _ F o l d e r 	 = " H a n d b � c k e r "  
  
 [ L i c e n s e A g r e e m e n t ]  
 T I T L E 	 = " L i c e n s a v t a l "  
 C B X _ A g r e e 	 = " J a g   g o d k � n n e r   v i l l k o r e n   i   a v t a l e t . "  
 I T M _ L a n g u a g e 	 = " S p r � k "  
 ; L N K _ P P 	 	 = " S e k r e t e s s p o l i c y "  
 ; U R L _ P P 	 	 = " h t t p : / / w w w . e p s o n . c o m / c g i - b i n / S t o r e / A b o u t P r i v a c y I n f o . j s p "  
 C O N F I R M 	 	 = " H a r   d u   l � s t   o c h   g o d k � n t   l i c e n s a v t a l e t   f � r   p r o g r a m v a r a n ? "  
  
 [ P r e p a r e ]  
 T I T L E 	 	 = " M a r k e r a   F � l j a n d e "  
 S U B _ T i t l e 	 = " "  
  
 [ S y s t e m C h e c k ]  
 T I T L E 	 = " K o n t r o l l e r a r   s y s t e m e t "  
 S U B _ T i t l e 	 = " "  
 T X T _ C h e c k P C 	 = " V � n t a   . . . "  
 T X T _ C h e c k N W 	 = " V � n t a   . . . "  
  
 ; �% 
 [ I n s t a l l O p t i o n ]  
 T I T L E 	 = " T i l l � g g s a v t a l "  
 S U B _ T i t l e 	 = " V � l j   v i l k a   i n s t a l l a t i o n s a l t e r n a t i v   d u   v i l l   a n v � n d a . "  
 T X T _ B o d y 	 = " "  
 C B X _ L a t e s t 	 = " L a d d a   n e r   d e n   s e n a s t e   p r o g r a m v a r a n   f r � n   E p s o n "  
 H L P _ L a t e s t 	 = " "  
 C B X _ S t a t u s 	 = " S t a t u s � v e r v a k n i n g   o c h   a u t o m a t i s k   u p p d a t e r a d   p r o g r a m v a r a   f r � n   E p s o n   % R E C O M M E N D E D % "  
 C B X _ G A 	 	 = " S k i c k a   a n v � n d n i n g s i n f o r m a t i o n   t i l l   E p s o n "  
 ; H L P _ G A 	 	 = " E p s o n   s a m l a r   i n   a n v � n d n i n g s i n f o r m a t i o n   f � r   a t t   f � r b � t t r a   p r o g r a m v a r a n s   k v a l i t e t   m e d   G o o g l e   A n a l y t i c s .   V i   s a m l a r   a l d r i g   i n   p e r s o n l i g   i n f o r m a t i o n . "  
 ; L N K _ G A 	 	 = " G o o g l e   A n a l y t i c s "  
 H L P _ G A 	 	 = " E p s o n   s a m l a r   i n   a n v � n d n i n g s i n f o r m a t i o n   f � r   a t t   f � r b � t t r a   k v a l i t e t e n   p �   v � r a   p r o d u k t e r   o c h   t j � n s t e r .   V i   s a m l a r   a l d r i g   i n   p e r s o n l i g   i n f o r m a t i o n . "  
 L N K _ G A 	 	 = " K l i c k a   h � r   f � r   m e r   u t f � r l i g   i n f o r m a t i o n "  
  
 [ I n s t a l l O p t i o n _ G A S u b ]  
 T I T L E 	 	 = " E p s o n   b e r   d i g   h j � l p a   o s s   m e d   a t t   f � r b � t t r a   v � r a   p r o d u k t e r   o c h   t j � n s t e r . "  
 C B X _ G A 	 	 = " T i l l � t   a t t   i n f o r m a t i o n   o m   p r o g r a m v a r u a n v � n d n i n g   s a m l a s   i n "  
 H L P _ G A 	 	 = " E p s o n   s a m l a r   i n   i n f o r m a t i o n   o m   p r o g r a m v a r u a n v � n d n i n g   m e d   G o o g l e   A n a l y t i c s . "  
 L N K _ G A 	 	 = " O m   G o o g l e   A n a l y t i c s "  
  
 C B X _ P L 	 	 = " T i l l � t   a t t   i n f o r m a t i o n   o m   p r o d u k t a n v � n d n i n g   s a m l a s   i n "  
 H L P _ P L 	 	 = " E p s o n   s a m l a r   i n   i n f o r m a t i o n   o m   p r o d u k t a n v � n d n i n g   m e d   p r o g r a m v a r a n   E p s o n   C u s t o m e r   R e s e a r c h . "  
 L N K _ P L 	 	 = " O m   p r o g r a m v a r a n   E p s o n   C u s t o m e r   R e s e a r c h "  
  
 C B X _ E R 	 	 = " E x p r e s s   P r o d u c t   R e g i s t r a t i o n "  
 H L P _ E R 	 	 = " E p s o n ' s   E x p r e s s   P r o d u c t   R e g i s t r a t i o n   p r o v i d e s   m a n y   v a l u a b l e   b e n e f i t s   t o   c u s t o m e r s ,   i n c l u d i n g   t e c h n i c a l   s u p p o r t   a n d   a d v i c e ,   f r e e   s o f t w a r e   u p d a t e s ,   e x c l u s i v e   o n l i n e   o f f e r s   a n d   n e w s   a b o u t   r e b a t e s ,   d i s c o u n t s ,   p r o d u c t   a n n o u n c e m e n t s   a n d   m o r e . "  
 L N K _ E R 	 	 = " A b o u t   E p s o n   E x p r e s s   P r o d u c t   R e g i s t r a t i o n "  
 T X T _ P P 	 	 = " B y   r e g i s t e r i n g   y o u r   p r o d u c t   y o u   a r e   p r o v i d i n g   y o u r   c o n s e n t   t o   E p s o n   A m e r i c a ,   I n c .   t o   u s e   y o u r   i n f o r m a t i o n   f o r   m a r k e t i n g   p u r p o s e s .   E p s o n   d o e s   n o t   s e l l   a n y   p e r s o n a l   i n f o r m a t i o n   t o   t h i r d   p a r t i e s .   Y o u   m a y   w i t h d r a w   y o u r   c o n s e n t   a t   a n y   t i m e .   V i e w   o u r   c o m p l e t e   < a   h r e f = " h t t p : / / w w w . e p s o n . c o m / c g i - b i n / S t o r e / A b o u t P r i v a c y I n f o . j s p " > p r i v a c y   p o l i c y < / a >   f o r   a d d i t i o n a l   i n f o r m a t i o n .   I f   y o u   a r e   a   C a l i f o r n i a   r e s i d e n t ,   p l e a s e   v i e w   o u r   < a   h r e f = " h t t p s : / / e p s o n . c o m / p r i v a c y - r i g h t s - c a l i f o r n i a " > C C P A   P r i v a c y   P o l i c y < / a > . "  
  
 [ I n s t a l l O p t i o n _ P L U R L ]  
 L N K _ U R L _ 1                     = " h t t p : / / s u p p o r t . e p s o n . n e t / P r i n t e r L o g g e r / s t 3 / i n d e x . p h p ? s e g = c p "  
 L N K _ U R L _ 2                     = " h t t p : / / s u p p o r t . e p s o n . n e t / P r i n t e r L o g g e r / s t 3 / i n d e x . p h p ? s e g = b p "  
 L N K _ U R L _ 3                     = " h t t p : / / s u p p o r t . e p s o n . n e t / P r i n t e r L o g g e r / s t 3 / i n d e x . p h p ? s e g = c p "  
 L N K _ U R L _ 4                     = " h t t p : / / s u p p o r t . e p s o n . n e t / P r i n t e r L o g g e r / s t 3 / i n d e x . p h p ? s e g = s c n "  
 L N K _ U R L _ 5                     = " h t t p : / / s u p p o r t . e p s o n . n e t / P r i n t e r L o g g e r / s t 3 / i n d e x . p h p ? s e g = l p "  
 L N K _ U R L _ 6                     = " h t t p : / / s u p p o r t . e p s o n . n e t / P r i n t e r L o g g e r / s t 3 / i n d e x . p h p ? s e g = s i d m "  
 L N K _ U R L _ 7                     = " h t t p : / / s u p p o r t . e p s o n . n e t / P r i n t e r L o g g e r / s t 3 / i n d e x . p h p ? s e g = l f p "  
  
 [ R e I n s t a l l ]  
 T I T L E 	 = " V � l j   T i l l v a l   a t t   i n s t a l l e r a "  
 S U B _ T i t l e 	 = " "  
 R B T _ E s s e n t i l a l   =   " I n s t a l l e r a   o m   d e n   p r o g r a m v a r a   s o m   k r � v s "  
 R B T _ A d d S o f t   =   " I n s t a l l e r a   v a l f r i   p r o g r a m v a r a "  
 R B T _ E x c h a n g e   = " K o n f i g u r e r a   d i n   p r o d u k t a n s l u t n i n g   i g e n \ n   ( i   h � n d e l s e   a v   n y   n � t v e r k s r o u t e r   e l l e r   b y t e   a v   U S B   t i l l   n � t v e r k   e l l e r   d y l i k t ) "  
  
 [ P r i n t e r L i s t ]  
 T I T L E 	 = " V � l j   v i l k e n   s o m   s k a   s t � l l a s   i n "  
 S U B _ T i t l e 	 = " "  
 R B T _ F i r s t 	 = " P r o d u k t   o c h   d a t o r "  
 H L P _ F i r s t 	 = " F � l j a n d e   s k � r m a r   v � g l e d e r   d i g   g e n o m   a t t   k o n f i g u r e r a   p r o d u k t e n   o c h   d a t o r n   f � r s t a   g � n g e n . "  
 R B T _ A d d i n g 	 = " E n d a s t   d a t o r n "  
 H L P _ A d d i n g 	 = " F � l j a n d e   p r o d u k t ( e r )   h a r   i d e n t i f i e r a t s   i   n � t v e r k e t .   V � l j   d e n   p r o d u k t   s o m   d u   v i l l   a n s l u t a   t i l l   o c h   k l i c k a   p �   % N E X T % .   O m   p r o d u k t e n   s o m   d u   v i l l   a n v � n d a   i n t e   v i s a s :   K o n t r o l l e r a   a t t   d e n   � r   p � s l a g e n   o c h   k l i c k a   p �   U p p d a t e r a . "  
 L S T _ M o d e l 	 = " P r o d u k t "  
 L S T _ M a c A d d r e s s 	 = " M A C - a d r e s s "  
 L S T _ I P A d d r e s s 	 = " I P - a d r e s s "  
 L N K _ I P _ M A N U A L 	 = " A v a n c e r a d   k o n f i g u r a t i o n "  
  
 [ I P M a n u a l S e t u p ]  
 T I T L E 	 = " L � g g   t i l l   s k r i v a r e   m e d   e n   s t a t i s k   I P - a d r e s s "  
 S U B _ T I T L E 	 = " "  
 T X T _ B o d y 	 = " A n g e   s k r i v a r e n s   I P - a d r e s s   n e d a n .   S e   t i l l   a t t   r e s e r v e r a   I P - a d r e s s e n   i   r o u t e r n s   i n s t � l l n i n g a r . "  
 I T M _ I P 	 = " I P - a d r e s s : "  
  
 [ H a r d w a r e S e t u p ]  
 T I T L E 	 = " I n s t a l l e r a "  
 S U B _ T i t l e 	 = " "  
  
 [ I n s t a l l E s s e n t i a l ]  
 T I T L E 	 = " I n s t a l l e r a   d e n   p r o g r a m v a r a   s o m   k r � v s "  
 T I T L E _ D L 	 = " H � m t a   d e n   p r o g r a m v a r a   s o m   k r � v s "  
 S U B _ T i t l e 	 = " "  
 T X T _ B o d y _ D L 	 = " L a d d a r   n e r   % s . . . "  
 T X T _ B o d y _ I N 	 = " I n s t a l l e r a r   % s . . . "  
 T X T _ B o d y _ U D 	 = " D e n   s e n a s t e   % s   � r   t i l l g � n g l i g . \ n V i l l   d u   i n s t a l l e r a ? "  
  
 [ F i r e w a l l G u i d e ]  
 T I T L E 	 	 = " K o n t r o l l e r a   d i n   s � k e r h e t s p r o g r a m v a r a "  
 T X T _ B o d y M a c 	 = " I f   y o u r   f i r e w a l l   s o f t w a r e   b l o c k s   t h e   n e t w o r k   c o n n e c t i o n   t o   t h e   p r o d u c t   o r   y o u   s e e   a   f i r e w a l l   a l e r t   s c r e e n ,   s e l e c t   t h e   o p t i o n   t h a t   a l l o w s   a c c e s s   t o   t h e   n e t w o r k   f o r   I n s t a l l   N a v i   i n   y o u r   f i r e w a l l   s o f t w a r e .   T h e n   c l i c k   [ % N E X T % ] . "  
  
 [ S e l e c t C o n n e c t ]  
 T I T L E 	 = " V � l j   d i n   a n s l u t n i n g s m e t o d "  
 S U B _ T i t l e 	 = " "  
 T X T _ B o d y 	 = " V � l j   h u r   d u   v i l l   a n s l u t a   p r o d u k t e n   t i l l   d i n   d a t o r ,   b � r b a r a   d a t o r   e l l e r   a n n a n   e n h e t . "  
 R B T _ W i f i 	 = " % W I F I % "  
 R B T _ W A C 	 = " % W I F I % "  
 R B T _ L A N 	 = " A n s l u t   v i a   t r � d b u n d e t   L A N   ( E t h e r n e t ) "  
 R B T _ U S B 	 = " A n s l u t   v i a   e n   U S B - k a b e l "  
  
 [ W i f i A u t o C o n n e c t ]  
 T I T L E 	 = " A n s l u t   t i l l   t r � d l � s t   L A N   a u t o m a t i s k t "  
  
 ; �% 
 [ W i f i A u t o C o n n e c t F P C ]  
 T I T L E _ N O 2 4 	 = " K u n d e   i n t e   h i t t a   d e n   t r � d l � s a   L A N - m i l j � n "  
  
 T I T L E _ S E T 2 4 	 = " V � l j   S S I D   o c h   l � s e n o r d   f � r   t r � d l � s t   L A N "  
 E X P _ S S I D 	 = " N � t v e r k s n a m n e t   ( S S I D )   a t t   s t � l l a   i n   f � r   p r o d u k t e n : "  
 E X P _ P W 	 	 = " L � s e n o r d : "  
 N O S S I D 	 	 = " V � l j   e t t   S S I D "  
  
 M S G _ S E T S S I D 	 = " A n s l u t   p r o d u k t e n   t i l l   S S I D   % s   i   d e n   t r � d l � s a   L A N - r o u t e r n . "  
 M S G _ S E T S S I D 2 	 = " V i l l   d u   a n s l u t a   p r o d u k t e n   a u t o m a t i s k t   t i l l   d e t t a   t r � d l � s a   L A N - S S I D :   [ % s ] "  
  
 M S G _ N O S E T 	 = " A n g e   l � s e n o r d e t . "  
 M S G _ E R R P W 	 = " L � s e n o r d e t   � r   o g i l t i g t .   A n g e   d e t   k o r r e k t a   v � r d e t . "  
 M S G _ E R R W A C 5 G 	 = " S S I D   e l l e r   l � s e n o r d   s o m   a n g i v i t s   f � r   p r o d u k t e n   k a n s k e   i n t e   � r   k o r r e k t . \ n K l i c k a   p �   [ % B A C K % ]   f � r   a t t   f � r s � k a   i g e n .   K l i c k a   p �   [ % N E X T % ]   f � r   a t t   k o n f i g u r e r a   m e d   e n   a n n a n   m e t o d . "  
  
 T I M E O U T _ C A U T I O N 	 = " O m   d e t   i n t r � f f a r   e t t   p r o d u k t f e l   s �   v � l j   A n s l u t   a u t o m a t i s k t   t i l l   W i - F i . "  
  
 [ W i f i A u t o C o n n e c t E r r o r ]  
 T I T L E 	 = " F e l   p �   t r � d l � s t   L A N - a n s l u t n i n g "  
 T I T L E _ W F D 	 = " F e l   p �   t r � d l � s t   L A N - a n s l u t n i n g "  
 S U B _ T i t l e 	 = " "  
 T X T _ B o d y 	 = " K u n d e   i n t e   a n s l u t a   t i l l   d i t t   n � t v e r k \ n K l i c k a   p �   [ % N E X T % ]   o c h   v � l j   e n   a n n a n   k o n f i g u r a t i o n s m e t o d   f � r   n � t v e r k e t . "  
 T X T _ B o d y A P 	 = " K u n d e   i n t e   a n s l u t a   t i l l   d i t t   n � t v e r k \ n K l i c k a   p �   [ % N E X T % ]   o c h   v � l j   e n   a n n a n   k o n f i g u r a t i o n s m e t o d   f � r   n � t v e r k e t . "  
 L N K _ V i d e o 	 = " W a t c h   V i d e o "  
  
 [ S S I D M a n u a l C o n n e c t ]  
 T I T L E 	 = " A n s l u t   t i l l   n � t v e r k   m a n u e l l t "  
 I T M _ S S I D 	 = " N � t v e r k s n a m n   ( S S I D ) : "  
 I T M _ P W 	 = " L � s e n o r d : "  
 B T N _ S h o w P W 	 = " V i s a   l � s e n o r d "  
 I T M _ P W E r r o r 	 = " I n t e   t i l l g � n g l i g "  
 I T M _ P W N o n e 	 = " O e t a b l e r a d "  
 L N K _ P u s h 	 = " I n s t a l l a t i o n   m e d   k n a p p t r y c k n i n g   f � r   W i - F i - n � t v e r k   ( W P S ) "  
 I T M _ S S I D _ P C 	 = " 5 G H z - n � t v e r k s n a m n   ( S S I D ) : "  
  
 [ E t h e r n e t C o n n e c t ]  
 T I T L E 	 = " A n s l u t   v i a   t r � d b u n d e t   L A N   ( E t h e r n e t ) "  
  
 [ U S B W i r e d C o n n e c t ]  
 T I T L E 	 = " A n s l u t   v i a   e n   U S B - k a b e l "  
 C B X _ L a t e r 	 = " A n s l u t   i n t e   n u "  
 G U I D E 	 = " I n s t a l l a t i o n e n   f o r t s � t t e r   a u t o m a t i s k t   n � r   e n   U S B - k a b e l   a n s l u t s . "  
  
 [ W i f i A u t o C o n n e c t W i t h U S B ]  
 T I T L E 	 = " A u t o m a t i s k   W i - F i - i n s t a l l a t i o n   ( t i l l f � l l i g   a n v � n d n i n g   a v   e n   U S B - k a b e l ) "  
 S U B _ T i t l e 	 = " "  
 C A U T I O N 	 = " K o p p l a   i n t e   u r   U S B - k a b e l n   f � r r � n   d u   o m b e d s   g � r a   d e t . "  
 G U I D E 	 = " I n s t a l l a t i o n e n   f o r t s � t t e r   a u t o m a t i s k t   n � r   e n   U S B - k a b e l   a n s l u t s . "  
  
 ; �% 
 [ U s e r S e l e c t C o n n e c t W r a p ]  
 T I T L E   = " V � l j   m e t o d   f � r   a t t   a n s l u t a   n � t v e r k e t "  
 S U B _ T i t l e 	 = " "  
 L N K _ P u s h 	 = " A n s l u t   m e d   W P S - k n a p p e n "  
 L N K _ W U S B 	 = " A n s l u t   m e d   t i l l f � l l i g   U S B - a n s l u t n i n g   ( h a   e n   U S B - k a b e l   t i l l   h a n d s ) "  
 L N K _ P a n e l 	 = " A n s l u t   g e n o m   a t t   a n g e   n � t v e r k s n a m n e t   ( S S I D )   o c h   l � s e n o r d e t   m a n u e l l t "  
 L N K _ I F S w i t c h 	 = " A n s l u t   g e n o m   a t t   a n g e   n � t v e r k s n a m n e t   ( S S I D )   o c h   l � s e n o r d e t   m a n u e l l t "  
  
 [ W i f i D i r e c t C o n n e c t ]  
 T I T L E 	 	 = " A n s l u t n i n g s i n s t � l l n i n g a r   f � r   W i - F i   D i r e c t   ( E n k e l   A P ) "  
 S U B _ T i t l e 	 = " "  
 T X T _ B o d y 	 = " D e t t a   u p p r � t t a r   e n   d i r e k t   W i - F i - a n s l u t n i n g   m e l l a n   d e n   h � r   d a t o r n   o c h   p r o d u k t e n . \ r \ n M e r   i n f o r m a t i o n   o m   W i - F i   D i r e c t   f i n n s   i   h a n d b o k e n . "  
  
 [ D i r e c t W i f i C o n n e c t ]  
 T I T L E 	 = " B e k r � f t a   a n s l u t n i n g s m e t o d e n "  
 S U B _ T i t l e 	 = " "  
 T X T _ B o d y 	 = " D e t t a   u p p r � t t a r   e n   d i r e k t   W i - F i - a n s l u t n i n g   m e l l a n   d e n   h � r   d a t o r n   o c h   p r o d u k t e n . \ r \ n M e r   i n f o r m a t i o n   o m   A P - l � g e   f i n n s   i   h a n d b o k e n . "  
  
 [ W F D M a n u a l ]  
 T I T L E 	 = " I n s t � l l n i n g   f � r   t r � d l � s   a n s l u t n i n g s h a n d b o k "  
 S U B _ T i t l e 	 = " "  
  
 [ P u s h B u t t o n C o n n e c t ]  
 T I T L E 	 = " A n s l u t   m e d   W P S - k n a p p e n "  
 T X T _ B o d y   = " A n s l u t   p r o d u k t e n   o c h   d e n   t r � d l � s a   r o u t e r n   a u t o m a t i s k t   g e n o m   a t t   t r y c k a   p �   d e n   t r � d l � s a   r o u t e r n s   k n a p p . "  
 S U B _ T i t l e 	 = " "  
 L N K _ A P m o d e 	 = " K l i c k a   h � r   o m   d i n   t r � d l � s a   r o u t e r   i n t e   s t � d e r   W P S - t r y c k k n a p p s f u n k t i o n e n "  
  
 [ A P m o d e M a n u a l S e t t i n g ]  
 T I T L E                 = " I n s t � l l n i n g   f � r   t r � d l � s   a n s l u t n i n g s h a n d b o k "  
  
 [ I P M a n u a l C o n n e c t ]  
 T I T L E 	 = " I n s t � l l n i n g   a v   n � t v e r k s p o r t "  
 S U B _ T i t l e 	 = " "  
 T X T _ S e t t i n g 	 = " S t � l l e r   i n   a n s l u t n i n g . . .   v � n t a . "  
  
 [ I n s t a l l N e t w o r k ]  
 T I T L E 	 = " L a d d a r   n e r   n � t v e r k s v e r k t y g "  
 S U B _ T i t l e 	 = " "  
 T X T _ B o d y _ D L 	 = " L a d d a r   n e r   % s . . . "  
 T X T _ B o d y _ I N 	 = " I n s t a l l e r a r   % s . . . "  
  
 ; �% 
 [ i f s _ i n p u t ]  
 T I T L E 	 	 = " A n s l u t   t i l l   n � t v e r k   m a n u e l l t "  
 T X T _ B o d y 	 = " "  
 I N P _ S S I D 	 = " S S I D   ( 2 , 4 G H z ) : "  
 I N P _ P W 	 	 = " L � s e n o r d : "  
 P L S _ S S I D 	 = " V � l j   e t t   S S I D "  
 P L S _ P W 	 	 = " W i - F i - n � t v e r k e t   % s   k r � v e r   e t t   l � s e n o r d . "  
 E R R _ T I T L E 	 = " F e l   p �   t r � d l � s t   L A N - a n s l u t n i n g "  
  
 [ N e t w o r k C o n n e c t e d ]  
 T I T L E 	 = " P r o d u k t   a n s l u t e n   t i l l   d i t t   n � t v e r k "  
 S U B _ T i t l e 	 = " "  
 S P I N F O 	 = " K o p p l a   u r   U S B - k a b e l n   o m   d u   h a r   a n v � n t   d e n   t i l l   n � t v e r k s i n s t a l l a t i o n e n . "  
 S P I N F O _ F U W 	 = " O b s :   L � t   U S B - k a b e l n   v a r a   a n s l u t e n   t i l l s   b a t t e r i e t   � r   f u l l a d d a t . "  
  
 [ L o c a l C o n n e c t e d ]  
 T I T L E 	 = " I n s t a l l a t i o n e n   � r   s l u t f � r d "  
 S U B _ T i t l e 	 = " "  
  
 ; �% 
 [ C o n n e c t e d G o E n d ]  
 T I T L E 2 	 	 = " O c h   n u . . . "  
 C K B _ E x p 1 	 = " P a r k o p p l a   s k a n n e r n   m e d   d a t o r n   f � r   a t t   s k a n n a   m e d   e n   k n a p p . "  
  
 ; �% 
 [ F W U p d a t e ]  
 T I T L E 	 	 = " K o n t r o l l e r a r   p r o g r a m v a r a n "  
 T I T L E 2 	 	 = " U p p d a t e r a r   p r o g r a m v a r a n "  
 T X T _ B o d y 	 = " V � n t a . . . S t � n g   i n t e   a v . "  
 T X T _ B o d y 2 	 = " V � n t a .   S t � n g   i n t e   a v   d i n   p r o d u k t   e l l e r   d a t o r .   P r o d u k t e n   k a n   s l u t a   f u n g e r a . "  
 E R R _ E S U 	 	 = " B � r j a r   k o n t r o l l e r a   d e n   i n b y g g d a   p r o g r a m v a r a n .   S t � n g   E p s o n   S o f t w a r e   U p d a t e r   o c h   k l i c k a   p �   [ O K ] . "  
 E R R _ V e r C h e c k 	 = " K u n d e   i n t e   k o n t r o l l e r a   d e n   i n b y g g d a   p r o g r a m v a r a n .   K o n t r o l l e r a   a t t   p r o d u k t e n   h a r   s l a g i t s   p �   o c h   a n s l u t i t s   t i l l   d a t o r n .   K l i c k a   s e d a n   p �   [ F � r s � k   i g e n ] .   K l i c k a   p �   [ H o p p a   � v e r ]   f � r   a t t   h o p p a   � v e r   i n s t � l l n i n g a r n a   f � r   P u s h   S c a n . "  
  
 ; �% 
 [ P a i r i n g ]  
 T I T L E 	 	 = " K o n f i g u r e r a   E n - k n a p p s s k a n n i n g "  
 T X T _ B o d y 	 = " V � n t a   . . . "  
 E R R _ A l r e a d y 	 = " S k a n n e r n   p a r k o p p l a s   m e d   e n   a n n a n   d a t o r .   V i l l   d u   p a r k o p p l a   s k a n n e r n   m e d   d e n   h � r   d a t o r n ? \ n E f t e r   p a r k o p p l i n g   k a n   d u   b � r j a   s k a n n a   g e n o m   a t t   t r y c k a   p �   s t a r t k n a p p e n   p �   s k a n n e r n   s �   s k i c k a s   d e t   d u   s k a n n a r   t i l l   d e n   d a t o r n . "  
  
 ; �% 
 [ F i r s t S c a n ]  
 T I T L E 	 	 = " T e s t a r   s k a n n i n g "  
  
 [ W a i t I n i t i a l C h a r g e ]  
 T I T L E 	 	 = " K o n t r o l l e r a   b l � c k i n i t i e r i n g s s t a t u s "  
 T X T _ B o d y 	 = " A n v � n d   i n t e   s k r i v a r e n   u n d e r   b l � c k i n i t i e r i n g e n .   V � n t a   t i l l s   p r o c e s s e n   � r   k l a r . "  
  
 [ T e s t P r i n t ]  
 T I T L E 	 = " S k r i v   u t   t e s t s i d a "  
 S U B _ T i t l e 	 = " "  
 L N K _ U t i l l i t y 	 = " F � r   p r o b l e m   m e d   u t s k r i f t s k v a l i t e t "  
 L N K _ L o t 4 	 = " I n f o r m a t i o n   o m   e f f e k t i v   e n e r g i f � r b r u k n i n g "  
 B T N _ P r i n t 	 = " S k r i v   u t   t e s t s i d a "  
  
 [ L o t 4 ]  
 T I T L E 	 = " I n f o r m a t i o n   o m   e f f e k t i v   e n e r g i f � r b r u k n i n g "  
 S U B _ T i t l e 	 = " "  
  
 [ I n v i t a t i o n ]  
 T I T L E 	 = " P r o d u k t r e g i s t r e r i n g   o n l i n e "  
 S U B _ T i t l e _ P R O D U C T 	 = " P r o d u k t n a m n "  
 S U B _ T i t l e _ S E R I A L 	 = " S e r i e n u m m e r "  
 R B T _ I n s t a l l 	 = " I n s t a l l e r a "  
 R B T _ D i s a g r e e 	 = " I n s t a l l e r a   i n t e "  
 R B T _ L a t e r 	 = " P � m i n n   m i g   s e n a r e "  
 T X T _ L o a d i n g 	 = " L a d d a r . . . "  
 T X T _ B o d y _ D L 	 = " H � m t a r   . . .   % s "  
 T X T _ B o d y _ I N 	 = " I n s t a l l e r a r   . . .   % s "  
 T X T _ R e g i o n 	 = " V � l j   d i t t   l a n d / r e g i o n . "  
 T X T _ N W _ E r r o r 	 = " K a n   i n t e   a n s l u t a   t i l l   i n t e r n e t .   K o n t r o l l e r a   d i n   a n s l u t n i n g   o c h   f � r s � k   i g e n . "  
  
 ; �% 
 [ F i n i s h ]  
 T I T L E 	 = " I n s t a l l a t i o n e n   � r   s l u t f � r d "  
 S U B _ T i t l e 	 = " "  
 T X T _ B o d y 	 = " D i n   p r o d u k t   � r   k l a r   a t t   a n v � n d a . "  
 T X T _ P M A 	 	 = " I f   y o u   e n r o l l e d   i n   a n   a u t o m a t i c   i n k   r e p l e n i s h m e n t   p r o g r a m ,   y o u   w i l l   c o n t i n u e   e n r o l l m e n t   a f t e r   y o u   e x i t   t h i s   i n s t a l l a t i o n   p r o g r a m . "  
 T I T L E 2 	 	 = " O c h   n u . . . "  
 C K B _ E x p 1 	 = " K o n t r o l l e r a   o m   d e t   f i n n s   u p p d a t e r a d   p r o g r a m v a r a "  
 C K B _ E x p 2 	 = " O n l i n e r e g i s t r e r i n g   f � r   d i n   p r o d u k t "  
  
 [ U n f i n i s h e d ]  
 T I T L E 	 = " I n s t a l l a t i o n e n   � r   k l a r "  
 S U B _ T i t l e 	 = " "  
 T X T _ B o d y 	 = " P r o g r a m v a r u i n s t a l l a t i o n e n   � r   k o m p l e t t . "  
  
 [ S e l e c t M o d e ]  
 T I T L E 	 	 = " H � m t a   W e b   I n s t a l l e r "  
 S U B _ T i t l e 	 = " V � l j   h u r   d u   v i l l   h � m t a   W e b   I n s t a l l e r . "  
 T X T _ B o d y 	 = " "  
 R B T _ W e b I n s t 	 = " I n s t a l l e r a   p �   d e n   h � r   d a t o r n "  
 H L P _ W e b I n s t 	 = " I n s t a l l e r a   n � d v � n d i g   p r o g r a m v a r a   o c h   a n s l u t   d e n n a   d a t o r . "  
 R B T _ S a v e F i l e 	 = " S p a r a   p �   e n   s � r s k i l d   p l a t s "  
 H L P _   S a v e F i l e 	 = " S p a r a   n � d v � n d i g   p r o g r a m v a r a   f � r   s e n a r e   i n s t a l l a t i o n   e l l e r   i n s t a l l e r a   p �   e n   d a t o r   s o m   i n t e   � r   a n s l u t e n   t i l l   i n t e r n e t . "  
 I T M _ S a v e i n 	 = " S p a r a   i "  
 I T M _   L a n g u a g e 	 = " S p r � k "  
  
 [ S a v e F i l e ]  
 T I T L E 	 	 = " S p a r a r   W e b   I n s t a l l e r "  
 S U B _ T i t l e 	 = " "  
 T X T _ B o d y 	 = " H � m t a r   . . .   % s "  
  
 [ S a v e F i n n i s h ]  
 T I T L E 	 	 = " W e b   I n s t a l l e r   h a r   s p a r a t s "  
 S U B _ T i t l e 	 = " "  
 T X T _ B o d y 	 = " W e b   I n s t a l l e r   h a r   s p a r a t s   t i l l   f � l j a n d e . "  
 I T M _ S a v e i n 	 = " F i l "  
 T X T _ R e a d 	 = " D u b b e l k l i c k a   p �   [ I n s t a l l N a v i . e x e ]   f � r   a t t   s t a r t a   i n s t a l l a t i o n e n . "  
  
 [ S y s t e m E r r o r ]  
 T I T L E 	 = " I n g e n   i n t e r n e t a n s l u t n i n g "  
 E R R _ A d m i n 	 = " D u   m � s t e   v a r a   i n l o g g a d   s o m   a d m i n i s t r a t � r   f � r   a t t   k u n n a   i n s t a l l e r a   p r o g r a m v a r a n . "  
 E R R _ O S 	 = " D i t t   o p e r a t i v s y s t e m   h a r   i n t e   s t � d   f � r   p r o g r a m v a r a n . "  
 E R R _ H D D 	 = " D e t   f i n n s   i n t e   t i l l r � c k l i g t   m e d   u t r y m m e   p �   d i t t   s y s t e m . \ r \ n V � l j   f � r r e   p r o g r a m   a t t   i n s t a l l e r a   e l l e r   f r i g � r   u t r y m m e   p �   d i t t   s y s t e m   o c h   i n s t a l l e r a   p r o g r a m m e n   i g e n . "  
  
 [ N W S e t t i n g E r r o r ]  
 T I T L E 	 = " N � t v e r k s k o n f i g u r a t i o n e n   a v b r � t s "  
 S U B _ T i t l e 	 = " S e   f e l s � k n i n g   n e d a n . "  
 T X T _ R e s t a r t 	 = " P r o d u k t n a m n e t   s o m   d u   v a l t   k a n   v a r a   f e l . "  
  
 [ T i m e O u t E r r o r ]  
 T I T L E 	 = " P r o d u k t e n   h i t t a d e s   i n t e "  
 S U B _ T i t l e 	 = " S e   f e l s � k n i n g   n e d a n . "  
 T X T _ R e s t a r t 	 = " P r o d u k t n a m n e t   s o m   d u   v a l t   k a n   v a r a   f e l . "  
  
 [ A b n o m a l E r r o r ]  
 T I T L E 	 = " F e l   v i d   a n s l u t n i n g   t i l l   n � t v e r k "  
 S U B _ T i t l e 	 = " S e   f e l s � k n i n g   n e d a n . "  
  
 [ W a i t C o n n e c t ]  
 T I T L E 	 = " N � t v e r k s k o n f i g u r a t i o n "  
 S U B _ T i t l e 	 = " H � m t a r   E p s o n N e t   S e t u p "  
 T X T _ B o d y 	 = " V � n t a   . . . "  
  
 [ W a i t S o f t w a r e ]  
 T I T L E 	 = " I n s t a l l e r a r   a p p l i k a t i o n s p r o g r a m v a r a "  
 S U B _ T i t l e 	 = " A n s l u t e r   t i l l   E p s o n   S o f t w a r e   U p d a t e r "  
 T X T _ B o d y 	 = " V � n t a   . . . "  
  
 [ N e t w o r k E r r o r ]  
 T I T L E 	 = " F e l   v i d   a n s l u t n i n g   t i l l   n � t v e r k "  
 S U B _ T i t l e 	 = " N � t v e r k e t s   g r � n s s n i t t   � r   i n t e   t i l l g � n g l i g t . "  
  
 [ W e b D o w n l o a d E r r o r ]  
 T I T L E 	 = " F e l   v i d   h � m t n i n g   a v   f i l "  
 E R R _ F a i l e d 	 = " K o n t r o l l e r a   I n t e r n e t a n s l u t n i n g e n   o c h   k l i c k a   O K .   K � r   s e d a n   i n s t a l l a t i o n s p r o g r a m m e t   i g e n . "  
 E R R _ R e t r y 	 = " K u n d e   i n t e   a n s l u t a   t i l l   I n t e r n e t .   V i l l   d u   f � r s � k a   i g e n ? "  
 E R R _ B u s y 	 = " K u n d e   i n t e   a n s l u t a   t i l l   s e r v e r n .   V i l l   d u   f � r s � k a   i g e n ? "  
 E R R _ C o m m 	 = " K o n t r o l l e r a   I n t e r n e t a n s l u t n i n g e n   o c h   k l i c k a   O K .   K � r   s e d a n   i n s t a l l a t i o n s p r o g r a m m e t   i g e n . "  
 B T N _ R E T R Y 	 = " F � r s � k   i g e n "  
  
 [ N W S e t t i n g C o m m o n ]  
 N O W _ S E T T I N G 	 = " I n s t a l l a t i o n   p � g � r .   V � n t a . . . "  
  
 [ N W S e t t i n g S t e p ]  
 S T E P I N F O _ B E G I N 	 = " S t a r t a   I n s t a l l a t i o n "  
 S T E P I N F O _ E U L A 	 = " L i c e n s a v t a l "  
 S T E P I N F O _ S Y S T E M C H E C K 	 = " S y s t e m k o n t r o l l "  
 S T E P I N F O _ I N S T A L L 	 = " I n s t a l l a t i o n "  
 S T E P I N F O _ C O N N E C T I O N 	 = " A n s l u t n i n g s i n s t � l l n i n g "  
 S T E P I N F O _ A D D I N S T A L L 	 = " K o m p l e t t e r a n d e   i n s t a l l a t i o n "  
 S T E P I N F O _ F I N I S H 	 = " S l u t f � r "  
 S T E P I N F O _ E N D 	 = " I n s t a l l a t i o n e n   � r   k l a r "  
  
 [ N W S e t t i n g B u t t o n ]  
 B U T T O N _ O K 	 = " O K "  
 B U T T O N _ C A N C E L 	 = " A v b r y t "  
 B U T T O N _ N E X T 	 = " N � s t a "  
 B U T T O N _ B A C K 	 = " B a k � t "  
 B U T T O N _ S K I P 	 = " H o p p a   � v e r "  
 T E X T _ Y E S 	 = " J a "  
 T E X T _ N O 	 	 = " N e j "  
  
 [ N W S e t t i n g W A C ]  
 T I T L E _ C S _ S I M P L E _ A P 	 = " P r o d u k t k o n f i g u r a t i o n   f � r   A n s l u t   a u t o m a t i s k t   t i l l   W i - F i "  
 S T E P 0 _ W A C 	 = " S � k e r   e f t e r   p r o d u k t . . . "  
 S T E P 1 _ W A C 	 = " K o n f i g u r e r a   n � t v e r k s i n f o r m a t i o n e n   f � r   p r o d u k t e n "  
 S T E P 2 _ W A C 	 = " K o n t r o l l e r a   a n s l u t n i n g e n "  
 S T E P 3 _ W A C 	 = " L � g g   t i l l   n � t v e r k s p r o d u k t e n   t i l l   d a t o r n "  
 S T E P 3 _ W A C _ M a c 	 = " � v r i g a   i n s t � l l n i n g a r "  
  
 [ N W S e t t i n g T C P I P ]  
 T I T L E _ T C P I P 	 = " I P - a d r e s s i n s t � l l n i n g a r "  
 L A B E L _ T C P I P 	 = " A k t u e l l   I P - a d r e s s   f � r   p r o d u k t e n   s t � l l s   i n   e n l i g t   n e d a n .   K l i c k a   p �   [ � n d r a ]   f � r   a t t   � n d r a   i n s t � l l n i n g a r n a   e l l e r   p �   [ N � s t a ]   f � r   a t t   f o r t s � t t a . "  
 L A B E L _ T C P I P _ S E T T I N G 	 = " I P - a d r e s s e n   f � r   p r o d u k t e n   � n d r a s   e n l i g t   h u r   d e t   v i s a s   h � r   n e d a n f � r .   K l i c k a   p �   [ N � s t a ]   f � r   a t t   f o r t s � t t a . \ n D u   k a n   � n g r a   � n d r i n g a r   g e n o m   a t t   k l i c k a   p �   [ � n g r a ] . "  
 R A D I O _ T C P I P _ A U T O 	 = " A u t o m a t i s k   k o n f i g u r e r i n g   a v   I P - a d r e s s   ( D H C P ) "  
 R A D I O _ T C P I P _ M A N U A L 	 = " M a n u e l l   k o n f i g u r e r i n g   a v   I P - a d r e s s   ( s t a t i s k   a d r e s s ) "  
 L A B E L _ T C P I P _ I P 	 = " I P - a d r e s s : "  
 L A B E L _ T C P I P _ S U B N E T 	 = " N � t m a s k : "  
 L A B E L _ T C P I P _ G A T E W A Y 	 = " S t a n d a r d g a t e w a y : "  
 B U T T O N _ T C P I P _ E D I T 	 = " � n d r a "  
 B U T T O N _ U N D O 	 = " � n g r a "  
 B U T T O N _ R E P R O B E 	 = " S � k   i g e n "  
  
 [ N W S e t t i n g T C P I P E r r o r ]  
 M S G _ I L L E G A L _ G A T E W A Y   =   " O g i l t i g   s t a n d a r d g a t e w a y . "  
 M S G _ I L L E G A L _ G A T E W A Y _ P A R E   =   " K o m b i n a t i o n e n   a v   s t a n d a r d g a t e w a y   o c h   n � t m a s k   � r   i n t e   g i l t i g . "  
 M S G _ I L L E G A L _ I P   =   " O g i l t i g   I P - a d r e s s . "  
 M S G _ I L L E G A L _ I P _ P A R E   =   " K o m b i n a t i o n e n   a v   I P - a d r e s s   o c h   n � t m a s k   � r   i n t e   g i l t i g . "  
 M S G _ I L L E G A L _ I P _ P A R E 2   =   " K o m b i n a t i o n e n   a v   I P - a d r e s s   o c h   s t a n d a r d g a t e w a y   � r   i n t e   g i l t i g . "  
 M S G _ I L L E G A L _ S U B N E T   =   " O g i l t i g   n � t m a s k . "  
  
 [ N W S e t t i n g T C P I P C o n f i r m ]  
 M S G _ Q U E S T I O N _ T C P I P _ S E T T I N G 	 = " K o n f i g u r a t i o n s m e t o d e n   e l l e r   I P - a d r e s s e n   f � r   p r o d u k t e n   � n d r a s . \ n F o r t s � t t a ? "  
  
 [ N W S e t t i n g S t o r a g e ]  
 T I T L E _ S T O R A G E _ A T T R I B U T E 	 = " F i l d e l n i n g s i n s t � l l n i n g a r "  
 L A B E L _ S T O R A G E 	 = " S t � l l   i n   s k r i v � t k o m s t   t i l l   e x t e r n a   l a g r i n g s e n h e t e r   s o m   e x e m p e l v i s   m i n n e s k o r t   e l l e r   U S B - m i n n e n   s o m   � r   a n s l u t n a   t i l l   p r o d u k t e n . \ n A n v � n d   i n t e   e x t e r n a   l a g r i n g s e n h e t e r   i n n a n   k o n f i g u r a t i o n e n   � r   s l u t f � r d .   D u   k a n   � n d r a   d e n   h � r   i n s t � l l n i n g e n   s e n a r e . "  
 T E X T _ R E A D W R I T E 	 = " W i - F i / n � t v e r k "  
 T E X T _ R E A D O N L Y 	 = " U S B "  
  
 [ N W S e t t i n g D r i v e r ]  
 T I T L E _ P R I N T S C A N 	 = " K o n f i g u r e r a   i n s t � l l n i n g a r "  
  
 [ N W S e t t i n g P r o d u c t S e a r c h ]  
 T I T L E _ P R O B E 	 = " S � k e r   e f t e r   p r o d u k t . . . "  
  
 [ N W S e t t i n g N o t F o u n d P r o d u c t s ]  
 M S G _ E R R O R _ N O _ P R I N T E R _ E A S Y M O D E 	 = " P r o d u k t e n   h i t t a d e s   i n t e .   K l i c k a   p �   [ O K ]   o c h   f � l j   i n s t r u k t i o n e r n a   p �   s k � r m e n   f � r   a t t   k � r a   k o n f i g u r a t i o n e n   i g e n . "  
  
 [ N W S e t t i n g S e l e c t M o d e l ]  
 T I T L E _ L I S T 	 = " V � l j   e n   p r o d u k t "  
 L A B E L _ L I S T 	 = " F � l j a n d e   p r o d u k t ( e r )   h a r   h i t t a t s   i   n � t v e r k e t .   V � l j   d e n   p r o d u k t   s o m   d u   v i l l   a n v � n d a   o c h   k l i c k a   p �   [ N � s t a ] .   O m   p r o d u k t e n   s o m   d u   v i l l   a n v � n d a   i n t e   v i s a s :   K o n t r o l l e r a   a t t   d e n   � r   p � s l a g e n . "  
 T E X T _ M O D E L 	 = " P r o d u k t n a m n "  
 T E X T _ S T A T U S 	 = " S t a t u s "  
 T E X T _ C O N N E C T S T Y L E 	 = " A n s l u t n i n g s t y p "  
 T E X T _ M A C 	 = " M A C - a d r e s s "  
 T E X T _ I P 	 = " I P - a d r e s s "  
 T E X T _ U S B 	 = " U S B "  
 T E X T _ W I R E D _ L A N 	 = " K a b e l a n s l u t e t   L A N "  
 T E X T _ W I R E L E S S _ L A N 	 = " T r � d l � s t   L A N "  
 T E X T _ S I M P L E _ A P 	 = " E n k e l   � t k o m s t p u n k t "  
  
 [ N W S e t t i n g U S B W A C ]  
 S T E P 0 _ U S B 	 = " A n g e   n � t v e r k s i n f o r m a t i o n "  
 S T E P 1 _ U S B 	 = " K o n f i g u r e r a   n � t v e r k s i n f o r m a t i o n e n   f � r   p r o d u k t e n "  
 S T E P 2 _ U S B 	 = " K o n t r o l l e r a   a n s l u t n i n g e n "  
 S T E P 3 _ U S B 	 = " L � g g   t i l l   n � t v e r k s p r o d u k t e n   t i l l   d a t o r n "  
 L A B E L _ L O C A L _ S E T T I N G S 	 = " D a t o r n   � r   a n s l u t e n   t i l l   f � l j a n d e   n � t v e r k   ( S S I D ) .   A n s l u t a   p r o d u k t e n   t i l l   n � t v e r k e t   ( S S I D ) ? "  
 L A B E L _ L O C A L _ S E T T I N G S _ S S I D 	 = " W i - F i - n � t v e r k s n a m n   ( S S I D ) : "  
 T I T L E _ S E N D I N G 	 = " S � n d e r   i n s t � l l n i n g a r "  
 T I T L E _ P O L L I N G 	 = " B e k r � f t a   a n s l u t n i n g e n "  
  
 [ N W S e t t i n g U S B W A C E r r o r ]  
 M S G _ E R R O R _ G E T D E T A I L 	 = " D e t   i n t r � f f a d e   e t t   f e l   v i d   k o m m u n i k a t i o n e n   m e d   p r o d u k t e n . \ n D e t   k a n   f i n n a s   e t t   p r o b l e m   m e d   p r o d u k t e n . \ n F � r s � k   a t t   s t � n g a   a v   p r o d u k t e n   o c h   s e d a n   s t a r t a   d e n   f � r   a t t   v � l j a   i n s t � l l n i n g a r n a   i g e n . "  
 M S G _ E R R O R _ C O N N E C T I N G _ 5 G H Z _ F R E Q U E N C Y _ B A N D 	 = " N � t v e r k s k a n a l e n   s o m   t i l l d e l a t s   t i l l   W i - F i - n � t v e r k   s t � d s   i n t e   a v   p r o d u k t e n .   D e t   k a n   i n a k t i v e r a   d i n   p r o d u k t s   W i - F i - a n s l u t n i n g . "  
  
 [ N W S e t t i n g A d m i n C o n f i r m ]  
 P A S S W D _ C A P T I O N 	 = " L � s e n o r d "  
 L A B E L _ P A S S W D 	 = " A n g e   a d m i n i s t r a t � r s l � s e n o r d e t   f � r   p r o d u k t e n . \ n O m   d u   i n t e   s t � l l t   i n   e t t   l � s e n o r d   a n g e r   d u   s e r i e n u m r e t   b a k i f r � n   a v   p r o d u k t e n . "  
 L A B E L _ P A S S W D 2 	 = " L � s e n o r d : "  
 T I T L E _ W I R E L E S S _ S E C U R I T Y _ A U T O 	 = " A n g e   a d m i n i s t r a t � r s l � s e n o r d "  
 M S G _ E R R O R _ S E T D E T A I L _ N O M A T C H _ P A S S W D 	 = " I n s t � l l n i n g e n   m i s s l y c k a d e s   e f t e r s o m   f e l   l � s e n o r d   a n g a v s . "  
 L A B E L _ P A S S W D _ N o C A 	 = " A n g e   a d m i n i s t r a t � r e n s   l � s e n o r d . "  
  
 [ B u t t o n T e x t ]  
 B T N _ Y e s                   = " J a "  
 B T N _ N o                     = " N e j "  
  
 [ N W H z E r r o r ]  
 M S G 	 	 = " A n s l u t n i n g e n   a v   p r o d u k t e n   m i s s l y c k a d e s   e f t e r s o m   d i n   d a t o r   � r   a n s l u t e n   t i l l   e t t   5 � G H z - S S I D   s o m   p r o d u k t e n   i n t e   h a r   s t � d   f � r .   A n s l u t   p r o d u k t e n   t i l l   e t t   2 , 4   G H z - S S I D   o c h   v � l j   s e d a n   p r o d u k t i n s t � l l n i n g a r n a . "  
  
 [ M a i n M a n u I t e m ]  
 T I T L E _ A B O U T _ A P P L I C A T I O N   =   " O m   % @ "  
 T I T L E _ H I D E _ A P P L I C A T I O N     =   " G � m   % @ "  
 T I T L E _ H I D E _ O T H E R S 	 	 =   " G � m   � v r i g a "  
 T I T L E _ S H O W _ A L L 	 	 	 =   " V i s a   a l l a "  
 T I T L E _ Q U I T _ A P P L I C A T I O N 	 =   " A v s l u t a   % @ "  
 T I T L E _ M I N I M I Z E 	 	 	 =   " M i n i m e r a "  
 T I T L E _ B R I N G _ A L L _ F R O N T 	 =   " L � g g   a l l a   � v e r s t "  
 T I T L E _ W I N D O W 	 =   " F � n s t e r "  
  
 [ S o f t w a r e U p d a t e ]  
 M A I N _ T I T L E 	 	 =   " I n s t a l l e r a r   v a l f r i   p r o g r a m v a r a "  
 S U B _ T i t l e 	 	 =   " "  
 C O L U M N _ T I T L E _ I N S T A L L 	 =   " I n s t a l l e r a "  
 C O L U M N _ T I T L E _ N A M E 	 	 =   " P r o g r a m "  
 C O L U M N _ T I T L E _ S T A T E 	 	 =   " S t a t u s "  
 C O L U M N _ T I T L E _ V E R S I O N 	 =   " V e r s i o n "  
 C O L U M N _ T I T L E _ S I Z E 	 	 =   " S t o r l e k "  
 S T A T E _ V A L U E _ N E W 	 	 	 =   " N y t t "  
 S T A T E _ V A L U E _ U P D A T E 	 	 =   " U p p d a t e r a "  
 S T A T E _ V A L U E _ I N S T A L L E D 	 =   " I n s t a l l e r a d "  
 B U T T O N _ N A M E _ I N S T A L L 	 	 =   " I n s t a l l e r a   % d   o b j e k t "  
 L A B E L _ T I T L E _ F R E E _ S P A C E 	 =   " L e d i g t   u t r y m m e   :   "  
 L A B E L _ T I T L E _ S U M 	 	 	 =   " T o t a l t   :   "  
 L A B E L _ T I T L E _ C H E C K 	 	 =   " K o n t r o l l e r a r   o m   d e t   f i n n s   p r o g r a m u p p d a t e r i n g a r . . . "  
 L A B E L _ T I T L E _ N O _ U P D A T E 	 =   " P r o g r a m v a r a n   � r   u p p d a t e r a d . "  
 L A B E L _ T I T L E _ R E Q U E S T 	 	 =   " A n s l u t e r   t i l l   s e r v e r . . . "  
 L A B E L _ T I T L E _ D O W N L O A D 	 =   " L a d d a r   n e r   % s . . . "  
 L A B E L _ T I T L E _ I N S T A L L 	 	 =   " I n s t a l l e r a r   % s . . . "  
 L A B E L _ U N I T _ M B 	 	 =   " G B "  
 L A B E L _ U N I T _ M B 	 	 =   " M B "  
  
 [ S o f t w a r e S e l e c t i o n ]  
 T I T L E 	 	 	 = " V � l j   P r o g r a m v a r a   a t t   i n s t a l l e r a "  
 C B X _ L a t e s t 	 	 = " L a d d a   n e r   d e n   s e n a s t e   p r o g r a m v a r a n   f r � n   E p s o n "  
 L A B E L _ T I T L E _ S U M 	 	 = " T o t a l t   :   "  
 L A B E L _ T I T L E _ F R E E _ S P A C E 	 = " L e d i g t   u t r y m m e   :   "  
 L A B E L _ T I T L E _ C H E C K 	 = " K o n t r o l l e r a r   o m   d e t   f i n n s   p r o g r a m u p p d a t e r i n g a r . . . "  
 L A B E L _ T I T L E _ N O _ U P D A T E 	 = " P r o g r a m v a r a n   � r   u p p d a t e r a d . "  
 L A B E L _ T I T L E _ R E Q U E S T 	 = " A n s l u t e r   t i l l   s e r v e r . . . "  
 L A B E L _ T I T L E _ D O W N L O A D 	 = " L a d d a r   n e r   % s . . . "  
 L A B E L _ T I T L E _ I N S T A L L 	 = " I n s t a l l e r a r   % s . . . "  
 L A B E L _ U N I T _ M B 	 	 = " M B "  
 L A B E L _ U N I T _ G B 	 	 = " G B "  
 L A B E L _ S T A T U S 	 	 = " S t a t u s   : "  
 L A B E L _ V E R S I O N 	 	 = " V e r s i o n   : "  
 L A B E L _ S I Z E 	 	 = " S t o r l e k   : "  
 S T A T U S _ N E W 	 	 = " N y t t "  
 S T A T U S _ U P D A T E 	 	 = " U p p d a t e r a "  
 S T A T U S _ I N S T A L L E D 	 = " I n s t a l l e r a d "  
 H L P _ B O T T O M _ L I S T 	 	 = " D u   k a n   i n t e   v � l j a   d e n   p r o g r a m v a r a   s o m   h a r   i n s t a l l e r a t s "  
 H L P _ B O T T O M _ L I S T 2 	 = " P r o g r a m v a r a   s o m   m a r k e r a t s   m e d   *   ( a s t e r i s k )   h a r   i n s t a l l e r a t s   o c h   k a n   i n t e   v � l j a s . "  
  
 [ C o n f i r m D r i v e r I n s t a l l ]  
 T X T _ B o d y   = " I n s t a l l e r a   e n   E P S O N - s k r i v a r d r i v r u t i n .   O m   d u   a n v � n d e r   e n   t r e d j e p a r t s d r i v r u t i n   k a n   d u   k l i c k a   p �   [ H o p p a   � v e r ] . "  
  
 [ e R e g _ W W ]  
 T I T L E 	 	 = " P r o d u k t r e g i s t r e r i n g   o n l i n e "  
 L S T _ R e g i o n 	 = " V � l j   d i t t   l a n d / r e g i o n . "  
 M S G _ M a i n 	 = " T a c k   f � r   a t t   d u   k � p t   e n   E p s o n - p r o d u k t .   V i   b e r   d i g   a t t   d u   r e g i s t r e r a r   E p s o n - p r o d u k t e n . \ r \ n V � l j   d i t t   l a n d / r e g i o n . "  
  
 [ C o n f i r m P u b l i c N e t w o r k ]  
 T X T _ B o d y 	 = " Y o u r   c o m p u t e r ' s   c u r r e n t   n e t w o r k   p r o f i l e   p r e v e n t s   d e v i c e   s h a r i n g .   T h i s   w i l l   d i s a b l e   s o m e   n e t w o r k   f u n c t i o n s   o n   y o u r   E p s o n   p r o d u c t ,   s u c h   a s   s c a n n i n g   f r o m   t h e   c o n t r o l   p a n e l .   F o r   a   n e t w o r k   y o u   t r u s t ,   i t   i s   r e c o m m e n d e d   t h a t   y o u   e n a b l e   s h a r i n g . \ n \ n W o u l d   y o u   l i k e   t o   e n a b l e   d e v i c e   s h a r i n g ? "  
  
 [ P r o d u c t R e g i s t r a t i o n ]  
 T I T L E   = " E x p r e s s   P r o d u c t   R e g i s t r a t i o n "  
 T I T L E _ E A I R E G   = " P r o d u k t r e g i s t r e r i n g "  
 T X T _ B o d y   = " C h e c k i n g   p r o d u c t   r e g i s t r a t i o n   s t a t u s . . . "  
 T X T _ B o d y _ P M A = " L a u n c h i n g   a u t o m a t i c   i n k   r e p l e n i s h m e n t   s e r v i c e   e n r o l l m e n t . . . "  
 T X T _ B o d y _ E A I R E G   = " S t a r t a r   p r o d u k t r e g i s t r e r i n g . . . "  
  
 [ R e s c u e M o d e ]  
 C O N F I R M 	 	 	 	 = " D e t   f i n n s   e t t   n y a r e   i n s t a l l a t i o n s p r o g r a m .   V i l l   d u   l a d d a   n e d   d e t ? "  
 M e s s a g e D o w n l o a d 	 	 = " D e t   n y a   i n s t a l l a t i o n s p r o g r a m m e t   l a d d a s   n e d .   V � n t a . . . \ n \ n I n s t a l l a t i o n s p r o g r a m m e t   b � r j a r   a u t o m a t i s k t   n � r   n e d l a d d n i n g e n   � r   s l u t f � r d . "  
 D o w n l o a d E r r o r 	 	 = " N e d l a d d n i n g e n   l y c k a d e s   i n t e .   V i l l   d u   f � r s � k a   i g e n ? "  
 